import PipeLineTypes::*;
import FIFO::*;
import FixedPoint::*;
import ClientServer::*;
import GetPut::*;
import Divide::*;

typedef struct {
    Frag a;
    Bool va;
    Frag b;
    Bool vb;
    Frag c;
    Bool vc;
    Frag d;
    Bool vd;
} FragWave deriving(Bits);

typedef Server#(
    Tuple2#(FragPos, FragPos),
    FragWave
) XiaoLinWu;


module mkFakeXiaoLinWu(XiaoLinWu);
	FIFO#(Tuple2#(FragPos, FragPos)) dummy <- mkFIFO;

	interface Put request;
		method Action put(Tuple2#(FragPos, FragPos) tup);
			dummy.enq(tup);
		endmethod
	endinterface
	
	interface Get response;
		method ActionValue#(FragWave) get();
			dummy.deq();
			Frag a = Frag{pos: tpl_1(dummy.first), intensity: maxBound};
			Frag b = Frag{pos: tpl_2(dummy.first), intensity: maxBound};
			return FragWave{a:a, va:True, b:b, vb:True, c:?, vc:False, d:?, vd:False};
		endmethod
	endinterface
endmodule

typedef struct {
	PixCoord x0;
	PixCoord x1;
	PixCoord y0;
	PixCoord y1;
	Fractional z0;
	Fractional z1;
	Bool swap;
} P2B deriving(Bits);

typedef struct {
	Fractional xdiff;
	Fractional ydiff;
	Fractional zdiff;
} P2A deriving(Bits);

typedef struct {
	Fractional k;
	Fractional k_inverse;
	Fractional kz;
	Fractional kz_alt;
} A2B deriving(Bits);

typedef struct {
	Fractional k;
} B2C deriving(Bits);

typedef struct {
	Fractional fky;
} C2D deriving(Bits);

typedef struct {
	FragPos l;
	FragPos r;
	Bool swaps;
} B2D deriving(Bits);

typedef struct {
	Bool xflip;
	Bool yflip;
} P2D deriving(Bits);

typedef struct {
	PixCoord x0;
	PixCoord y0;
	Fractional z0;
	PixCoord x1;
	PixCoord y1;
	Fractional z1;
	Fractional kz;
} B2R deriving(Bits);

typedef struct {
	Offset ky;
	Offset oD;
	Bool xflip;
	Bool yflip;
	Bool swaps;
} D2R deriving(Bits);

module mkXiaoLinWu(XiaoLinWu);

    FIFO#(FragWave) outFIFO <- mkFIFO;
    
    FIFO#(P2A) p2aFIFO <- mkFIFO;
    FIFO#(A2B) a2bFIFO <- mkFIFO;
    FIFO#(P2B) p2bFIFO <- mkFIFO;
    FIFO#(B2C) b2cFIFO <- mkFIFO;
    FIFO#(P2D) p2dFIFO <- mkFIFO;
    FIFO#(C2D) c2dFIFO <- mkFIFO;
    FIFO#(B2D) b2dFIFO <- mkFIFO;
    
    // These are the values generated by the initialization phase,
    // and used by the interpolation phase
    FIFO#(B2R) b2rFIFO <- mkFIFO;
    FIFO#(D2R) d2rFIFO <- mkFIFO;
    
    // State used by the interpolation stage
    Reg#(Bool) is_interpolating <- mkReg(False);
    Reg#(PixCoord) x0 <- mkRegU;
    Reg#(PixCoord) y0 <- mkRegU;
    Reg#(Fractional) z0 <- mkRegU;
    Reg#(PixCoord) x1 <- mkRegU;
    Reg#(PixCoord) y1 <- mkRegU;
    Reg#(Fractional) z1 <- mkRegU;
    Reg#(Fractional) kz <- mkRegU;
    Reg#(Offset) ky <- mkRegU;
    Reg#(Offset) oD <- mkRegU;
    Reg#(Offset) prev_oD <- mkRegU;
    
    Reg#(Bool) xflip <- mkRegU;
    Reg#(Bool) yflip <- mkRegU;
    Reg#(Bool) swaps <- mkRegU;
    
    Server#(Tuple2#(Int#(32),Int#(16)), Tuple2#(Int#(16),Int#(16))) d1 <- mkSignedDivider(1);
    Server#(Tuple2#(Int#(32),Int#(16)), Tuple2#(Int#(16),Int#(16))) d2 <- mkSignedDivider(1);
    Server#(Tuple2#(Int#(32),Int#(16)), Tuple2#(Int#(16),Int#(16))) d3 <- mkSignedDivider(1);
    Server#(Tuple2#(Int#(32),Int#(16)), Tuple2#(Int#(16),Int#(16))) d4 <- mkSignedDivider(1);
    
    function Tuple2#(FragPos, FragPos) descramble(FragPos a, FragPos b,
    											  Bool xf, Bool yf, Bool sw);
        PixCoord tx0 = (sw) ? a.y : a.x;
        PixCoord ty0 = (sw) ? a.x : a.y;
        PixCoord tx1 = (sw) ? b.y : b.x;
        PixCoord ty1 = (sw) ? b.x : b.y;
        PixCoord oy1 = (yf) ? ty0 : ty1;
        PixCoord oy0 = (yf) ? ty1 : ty0;
        PixCoord ox1 = (xf) ? tx0 : tx1;
        PixCoord ox0 = (xf) ? tx1 : tx0;
        return tuple2(FragPos{x:ox0, y:oy0, z:a.z},
                      FragPos{x:ox1, y:oy1, z:b.z});
    endfunction

	// interpolation state
	rule begin_interpolate(!is_interpolating);
		let b2r = b2rFIFO.first();
		let d2r = d2rFIFO.first();
		b2rFIFO.deq();
		d2rFIFO.deq();
		
		is_interpolating <= True;

		y0 <= b2r.y0;
		y1 <= b2r.y1;
		kz <= b2r.kz;
		ky <= d2r.ky;
		prev_oD <= d2r.oD;
		xflip <= d2r.xflip;
		yflip <= d2r.yflip;
		swaps <= d2r.swaps;
		
		oD <= d2r.oD + d2r.ky;
		x0 <= b2r.x0 + 1;
		x1 <= b2r.x1 - 1;
		z0 <= b2r.z0 + b2r.kz;
		z1 <= b2r.z1 - b2r.kz;
	endrule
	
	rule interpolate(is_interpolating);
		let thisy0 = y0;
		let thisy1 = y1;
		if ((oD <= prev_oD) && ky != 0) begin
			thisy0 = thisy0 + 1;
			thisy1 = thisy1 - 1;
		end
		
		// Intensity is calculated from the current offset value (oD)
		Intensity intensity = truncate(oD >> (valueOf(N_BITS) - valueOf(M_BITS)) );
        Intensity invertedI = ~intensity;
        
        // Left, right, up, down fragments (up is above left, down is below right)
        FragPos l = FragPos{x:x0, y:thisy0, z:z0};
        FragPos r = FragPos{x:x1, y:thisy1, z:z1};
        FragPos u = FragPos{x:x0, y:thisy0+1, z:z0};
        FragPos d = FragPos{x:x1, y:thisy1-1, z:z1};
        
        let outp = descramble(l, r, xflip, yflip, swaps);
        let outs = descramble(u, d, xflip, yflip, swaps);
        
        // Enqueue wave of Fragments
        FragWave outwave;
        outwave.a = Frag{pos: tpl_1(outp), intensity: invertedI};
        outwave.va = True;
        outwave.b = Frag{pos: tpl_2(outp), intensity: invertedI};
        outwave.vb = True;
        outwave.c = Frag{pos: tpl_1(outs), intensity: intensity};
        outwave.vc = True;
        outwave.d = Frag{pos: tpl_2(outs), intensity: intensity};
        outwave.vd = True;
        
        if (x0 > x1) begin
        	is_interpolating <= False;
        end else begin
        	outFIFO.enq(outwave);
        end
        // Following logically in else block but in that case
        // is inconsequential anyway
        prev_oD <= oD;
        oD <= oD + ky;
		x0 <= x0 + 1;
		x1 <= x1 - 1;
		y0 <= thisy0;
		y1 <= thisy1;
		z0 <= z0 + kz;
		z1 <= z1 - kz;
	endrule
    
    rule a_to_div;
    	// get input fifo
    	let p = p2aFIFO.first();
    	// dequeue input fifo
		p2aFIFO.deq();
		
		// enqueue division
		Int#(16) x_small = unpack({p.xdiff.i,p.xdiff.f});
		Int#(16) y_small = unpack({p.ydiff.i,p.ydiff.f});
		Int#(24) x_medium = unpack({pack(x_small),0});
		Int#(24) y_medium = unpack({pack(y_small),0});
		Int#(24) z_medium = unpack({p.zdiff.i,p.zdiff.f,0});
		Int#(32) x_big = extend(x_medium);
		Int#(32) y_big = extend(y_medium);
		Int#(32) z_big = extend(z_medium);
		d1.request.put(tuple2(y_big,x_small));
		d2.request.put(tuple2(x_big,y_small));
		d3.request.put(tuple2(z_big,x_small));
		d4.request.put(tuple2(z_big,y_small));
    endrule
    
    rule div_to_b;
    	let r1 <- d1.response.get();
    	let r2 <- d2.response.get();
    	let r3 <- d3.response.get();
    	let r4 <- d4.response.get();
    	let p1 = pack(tpl_1(r1));
    	let p2 = pack(tpl_1(r2));
    	let p3 = pack(tpl_1(r3));
    	let p4 = pack(tpl_1(r4));
    	let k 		 = Fractional{i:p1[15:8],f:p1[7:0]};
    	let inverseK = Fractional{i:p2[15:8],f:p2[7:0]};
    	let k_z 	 = Fractional{i:p3[15:8],f:p3[7:0]};
    	let k_z_alt  = Fractional{i:p4[15:8],f:p4[7:0]};
    	a2bFIFO.enq(A2B{k:k,k_inverse:inverseK,kz:k_z,kz_alt:k_z_alt});
    endrule
    
    rule b;
    	// Get input fifos
    	let a2b = a2bFIFO.first();
    	let p2b = p2bFIFO.first();
    	// deque input fifos
    	a2bFIFO.deq();
		p2bFIFO.deq();
    	
		//let thisSwaps = (a2b.k > 1.0);
		let thisSwaps = p2b.swap;
		let thisx0 = (thisSwaps) ? p2b.y0 : p2b.x0;
		let thisx1 = (thisSwaps) ? p2b.y1 : p2b.x1;
		let thisy0 = (thisSwaps) ? p2b.x0 : p2b.y0;
		let thisy1 = (thisSwaps) ? p2b.x1 : p2b.y1;
		let thisz0 = (thisSwaps) ? p2b.z1 : p2b.z0;
		let thisz1 = (thisSwaps) ? p2b.z0 : p2b.z1;
		
		let thisk = (thisSwaps) ? a2b.k_inverse : a2b.k;
		let thiskz = (thisSwaps) ? a2b.kz_alt : a2b.kz;
		
		// Left, right endpoints
		FragPos l = FragPos{x:thisx0, y:thisy0, z:thisz0};
		FragPos r = FragPos{x:thisx1, y:thisy1, z:thisz1};
		
		// enqueue output fifos
		b2dFIFO.enq(B2D{l:l,r:r,swaps:thisSwaps});
		b2cFIFO.enq(B2C{k:thisk});
		// enqueue to interpolation stage
		b2rFIFO.enq(B2R{x0:thisx0,y0:thisy0,z0:thisz0,
						x1:thisx1,y1:thisy1,z1:thisz1});
    endrule
    
    rule c;
    	// get input fifo
    	let b2c = b2cFIFO.first();
    	// dequeue input fifo
    	b2cFIFO.deq();
    	
    	Offset maxval = maxBound;
    	Fractional fmaxval = Fractional{i:{'0, pack(maxval)[13:7]}, f:{pack(maxval)[6:0], '0}};
    	Fractional fractky = b2c.k * fmaxval;
    	
    	// enqueue output fifo
    	c2dFIFO.enq(C2D{fky:fractky});
    endrule
    
    rule d;
    	// get input fifos
    	let p2d = p2dFIFO.first();
    	let b2d = b2dFIFO.first();
    	let c2d = c2dFIFO.first();
    	// dequeue input fifos
    	p2dFIFO.deq();
    	b2dFIFO.deq();
    	c2dFIFO.deq();
    	
    	let in_xflip = p2d.xflip;
    	let in_yflip = p2d.yflip;
    	let in_swaps = b2d.swaps;
    	let outs = descramble(b2d.l, b2d.r,
    						  in_xflip, in_yflip, in_swaps);

		// Make a new FragWave and build it
		FragWave outwave;
		outwave.a = Frag{pos: tpl_1(outs), intensity: maxBound};
		outwave.va = True;
		outwave.b = Frag{pos: tpl_2(outs), intensity: maxBound};
		outwave.vb = True;
		outwave.c = ?;
		outwave.vc = False;
		outwave.d = ?;
		outwave.vd = False;
		outFIFO.enq(outwave);
			
		Offset thisky = unpack({c2d.fky.i[6:0], c2d.fky.f[7:1]});
		
		// enqueue to interpolation stage
		d2rFIFO.enq(D2R{ky:thisky,oD:0,xflip:in_xflip,yflip:in_yflip,swaps:in_swaps});
    endrule

	interface Put request;
	    method Action put(Tuple2#(FragPos, FragPos) tup);
	    	let a = tpl_1(tup); // pipeline
	    	let b = tpl_2(tup); // pipeline
			let xf = (a.x > b.x);
			let yf = (a.y > b.y);
	
			let tx0 = (xf) ? b.x : a.x; // pipeline
			let tx1 = (xf) ? a.x : b.x; // pipeline
			let ty0 = (yf) ? b.y : a.y; // pipeline
			let ty1 = (yf) ? a.y : b.y; // pipeline

			// Subtraction
			Bit#(10) xdiff_ten = extend(pack(tx1)) - extend(pack(tx0));
			Bit#(10) ydiff_ten = extend(pack(ty1)) - extend(pack(ty0));
			// Just wires
			Bit#(8) xdiff_integer = {'0, xdiff_ten[9:3]};
			Bit#(8) xdiff_fraction = {xdiff_ten[2:0], '0};
			Bit#(8) ydiff_integer = {'0, ydiff_ten[9:3]};
			Bit#(8) ydiff_fraction = {ydiff_ten[2:0], '0};
			Fractional xdiff = Fractional{i:xdiff_integer, f:xdiff_fraction}; // pipeline
			Fractional ydiff = Fractional{i:ydiff_integer, f:ydiff_fraction}; // pipeline
			Fractional zdiff = b.z - a.z; // pipeline
			
			//test
			Bool mSwaps = ydiff > xdiff;
			
			// Give data to next steps of line initialization
			p2bFIFO.enq(P2B{x0:tx0,x1:tx1,y0:ty0,y1:ty1,z0:a.z,z1:b.z,swap:mSwaps});
			p2aFIFO.enq(P2A{xdiff:xdiff,ydiff:ydiff,zdiff:zdiff});
			p2dFIFO.enq(P2D{xflip:xf, yflip:yf});
	    endmethod
	endinterface
	
    interface response = toGet(outFIFO);
endmodule


/*
		$display("HW: XiaoLinWu: line started, outwave enqueued");
		
		$display("tx0: %d, ty0: %d, tx1: %d, ty1: %d", tx0, ty0, tx1, ty1);
		$display("ixdiff: %d", ixdiff);
		$write("xdiff: "); fxptWrite(3, xdiff*32); $display(" ");
		$write("ydiff: "); fxptWrite(3, ydiff*32); $display(" ");
		$write("k: "); fxptWrite(3, k); $display(" ");
		$write("fractky: "); fxptWrite(3, fractky); $display(" ");
		$write("fractMaxVal: "); fxptWrite(3, fractMaxVal); $display(" ");
		$display("fractky.i: %b", fractky.i);
		$display("fractky.i[5:0]: %b", fractky.i[5:0]);
		$display("ky: %d", thisky);
		$display("maxval: %d", maxval);
		*/
